// fir.v

// Generated using ACDS version 22.1 915

`timescale 1 ps / 1 ps
module fir (
		input  wire [5:0]   coeff_in_address, //         avalon_mm_slave.address
		input  wire         coeff_in_read,    //                        .read
		output wire [0:0]   coeff_out_valid,  //                        .readdatavalid
		output wire [15:0]  coeff_out_data,   //                        .readdata
		input  wire [0:0]   coeff_in_we,      //                        .write
		input  wire [15:0]  coeff_in_data,    //                        .writedata
		input  wire [79:0]  ast_sink_data,    //   avalon_streaming_sink.data
		input  wire         ast_sink_valid,   //                        .valid
		input  wire [1:0]   ast_sink_error,   //                        .error
		output wire [219:0] ast_source_data,  // avalon_streaming_source.data
		output wire         ast_source_valid, //                        .valid
		output wire [1:0]   ast_source_error, //                        .error
		input  wire         clk,              //                     clk.clk
		input  wire         coeff_in_clk,     //             coeff_clock.clk
		input  wire         coeff_in_areset,  //             coeff_reset.reset_n
		input  wire         reset_n           //                     rst.reset_n
	);

	fir_fir_compiler_ii_0 fir_compiler_ii_0 (
		.clk              (clk),              //                     clk.clk
		.reset_n          (reset_n),          //                     rst.reset_n
		.ast_sink_data    (ast_sink_data),    //   avalon_streaming_sink.data
		.ast_sink_valid   (ast_sink_valid),   //                        .valid
		.ast_sink_error   (ast_sink_error),   //                        .error
		.ast_source_data  (ast_source_data),  // avalon_streaming_source.data
		.ast_source_valid (ast_source_valid), //                        .valid
		.ast_source_error (ast_source_error), //                        .error
		.coeff_in_clk     (coeff_in_clk),     //             coeff_clock.clk
		.coeff_in_areset  (coeff_in_areset),  //             coeff_reset.reset_n
		.coeff_in_address (coeff_in_address), //         avalon_mm_slave.address
		.coeff_in_read    (coeff_in_read),    //                        .read
		.coeff_out_valid  (coeff_out_valid),  //                        .readdatavalid
		.coeff_out_data   (coeff_out_data),   //                        .readdata
		.coeff_in_we      (coeff_in_we),      //                        .write
		.coeff_in_data    (coeff_in_data)     //                        .writedata
	);

endmodule
